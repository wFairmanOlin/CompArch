// Simple Verilog Test
module hello_test ();
initial begin
	$display("Hellow, Comparch!");
end
endmodule
